aottaviano@maipo.ee.ethz.ch.22822:1604756657